`timescale 1ns/1ns

module Sumador4(
    input [31:0]sum_in1,
    output [31:0]suma_out
);

assign suma_out=sum_in1+4;

endmodule
